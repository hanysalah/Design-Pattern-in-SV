class ParentClass;

   virtual function ParentClass clone();
   endfunction // clone

endclass // ParentClass
