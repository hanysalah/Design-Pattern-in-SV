package non_touch_package;

`include "parent.sv"
`include "childClasses.sv"
`include "childChildClasses.sv"

endpackage