virtual class StrategyObjectClass;
endclass


class StrategyObjectOneClass extends StrategyObjectClass;
endclass


class StrategyObjectTwoClass extends StrategyObjectClass;
endclass