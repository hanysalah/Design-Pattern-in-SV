class child1Child1 extends child1;

endclass

class child2Child1 extends child1;

endclass

class child1Child2 extends child2;

endclass

class child2Child2 extends child2;

endclass