class child2_extension extends child2;

  virtual function void do_FuncVirtual();
    $display("Here is the extended implementation in Child 2");
  endfunction

endclass